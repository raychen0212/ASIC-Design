mg35@ecegrid-thin5.ecn.purdue.edu.46123:1608406941