// $Id: $
// File name:   tb_apb_uart_rx.sv
// Created:     3/22/2021
// Author:      Jhen-Ruei Chen
// Lab Section: 337-08
// Version:     1.0  Initial Design Entry
// Description: Test bench for apb UART
